module projetorelogio (input a, output o);

	

endmodule
